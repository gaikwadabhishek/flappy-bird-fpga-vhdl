library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.MY.all;

ENTITY SYNC IS
PORT (
	CLK: IN STD_LOGIC;
	HSYNC, VSYNC: OUT STD_LOGIC;
	R, G, B : OUT STD_LOGIC_VECTOR(3 downto 0);
	KEYS: IN STD_LOGIC_VECTOR(3 downto 0);
	S: IN STD_LOGIC_VECTOR(1 downto 0)
);
END SYNC;

ARCHITECTURE MAIN OF SYNC IS
SIGNAL RGB: STD_LOGIC_VECTOR(3 downto 0);
SIGNAL DRAW1, DRAW2, DRAW3, DRAW4, DRAW5, DRAW6, DRAW7, DRAW8, DRAW9, DRAW10, DRAW11, DRAW12, DRAW13: STD_LOGIC;
SIGNAL START, STOP: STD_LOGIC := '0';
SIGNAL SQ_X1, SQ_Y1: INTEGER RANGE 0 TO 1688:=600;
SIGNAL SQ_X2, SQ_Y2: INTEGER RANGE 0 TO 1688:=800;

SIGNAL PB_X1, PA_X1: INTEGER RANGE 0 TO 1688:=0;
SIGNAL PA_Y1: INTEGER RANGE 0 TO 1688:=0;
SIGNAL PB_Y1: INTEGER RANGE 0 TO 1688:=1688;

SIGNAL PB_X2, PA_X2: INTEGER RANGE 0 TO 1688:=408;
SIGNAL PA_Y2: INTEGER RANGE 0 TO 1688:=000;
SIGNAL PB_Y2: INTEGER RANGE 0 TO 1688:=1688;

SIGNAL PB_X3, PA_X3: INTEGER RANGE 0 TO 1688:=808;
SIGNAL PA_Y3: INTEGER RANGE 0 TO 1688:=000;
SIGNAL PB_Y3: INTEGER RANGE 0 TO 1688:=1688;

SIGNAL PB_X4, PA_X4: INTEGER RANGE 0 TO 1688:=1208;
SIGNAL PA_Y4: INTEGER RANGE 0 TO 1688:=000;
SIGNAL PB_Y4: INTEGER RANGE 0 TO 1688:=1688;

SIGNAL PB_X5, PA_X5: INTEGER RANGE 0 TO 1688:=1688;
SIGNAL PA_Y5: INTEGER RANGE 0 TO 1688:=000;
SIGNAL PB_Y5: INTEGER RANGE 0 TO 1688:=1688;

SIGNAL PB_X6, PA_X6: INTEGER RANGE 0 TO 1688:=1688;
SIGNAL PA_Y6: INTEGER RANGE 0 TO 1688:=000;
SIGNAL PB_Y6: INTEGER RANGE 0 TO 1688:=1688;

SIGNAL HPOS: INTEGER RANGE 0 TO 1688:=0;
SIGNAL VPOS: INTEGER RANGE 0 TO 1066:=0;
BEGIN
SQ(HPOS, VPOS, SQ_X1, SQ_Y1, RGB, DRAW1);
PIPE_BELOW(HPOS, VPOS, PB_X1, PB_Y1, RGB, DRAW2);
PIPE_ABOVE(HPOS, VPOS, PA_X1, PA_Y1, RGB, DRAW3);

PIPE_BELOW(HPOS, VPOS, PB_X2, PB_Y2, RGB, DRAW4);
PIPE_ABOVE(HPOS, VPOS, PA_X2, PA_Y2, RGB, DRAW5);

PIPE_BELOW(HPOS, VPOS, PB_X3, PB_Y3, RGB, DRAW6);
PIPE_ABOVE(HPOS, VPOS, PA_X3, PA_Y3, RGB, DRAW7);

PIPE_BELOW(HPOS, VPOS, PB_X4, PB_Y4, RGB, DRAW8);
PIPE_ABOVE(HPOS, VPOS, PA_X4, PA_Y4, RGB, DRAW9);

PIPE_BELOW(HPOS, VPOS, PB_X5, PB_Y5, RGB, DRAW10);
PIPE_ABOVE(HPOS, VPOS, PA_X5, PA_Y5, RGB, DRAW11);

PIPE_BELOW(HPOS, VPOS, PB_X6, PB_Y6, RGB, DRAW12);
PIPE_ABOVE(HPOS, VPOS, PA_X6, PA_Y6, RGB, DRAW13);


PROCESS (CLK)
BEGIN
IF (CLK'EVENT AND CLK='1') THEN

	IF (DRAW1='1') THEN
		R <= (OTHERS => '1');
		G <= (OTHERS => '1');
		B <= (OTHERS => '1');
	END IF;

	IF PB_X1 < 10 THEN
		PA_Y1 <= 650;
		PB_Y1 <= PA_Y1 + 275;
	END IF;
	
	IF PB_X2 < 10 THEN
		PA_Y2 <= 350;
		PB_Y2 <= PA_Y2 + 275;
	END IF;
	
	IF PB_X3 < 10 THEN
		PA_Y3 <= 500;
		PB_Y3 <= PA_Y3 + 275;
	END IF;
	
	IF PB_X4 < 10 THEN
		PA_Y4 <= 200;
		PB_Y4 <= PA_Y4 + 275;
	END IF;
	
	IF PB_X5 < 10 THEN
		PA_Y5 <=650;
		PB_Y5 <= PA_Y5 + 275;
	END IF;
	
	IF (DRAW2='1' OR DRAW3='1' OR DRAW4='1' OR DRAW5='1' OR DRAW6='1' OR DRAW7='1' OR DRAW8='1'OR DRAW9='1' OR DRAW10='1' OR DRAW11='1' OR DRAW12='1' OR DRAW13='1') THEN
			R <= (OTHERS => '0');
			G <= (OTHERS => '1');
			B <= (OTHERS => '0');
	END IF;
	
	IF (DRAW1 = '0' AND DRAW2 = '0' AND DRAW3 = '0' AND DRAW4 = '0' AND DRAW5 = '0' AND DRAW6 = '0' AND DRAW7 = '0' AND DRAW7 = '0' AND DRAW8 = '0' AND DRAW9 = '0' AND DRAW10 = '0' AND DRAW11 = '0' AND DRAW12 = '0' AND DRAW13 = '0') THEN
		R <= (OTHERS => '0');
		G <= (OTHERS => '0');
		B <= (OTHERS => '1');
	END IF;
	
	IF (DRAW1 = '1' AND (DRAW2='1' OR DRAW3='1' OR DRAW4='1' OR DRAW5='1' OR DRAW6='1' OR DRAW7='1' OR DRAW8='1'OR DRAW9='1' OR DRAW10='1' OR DRAW11='1' OR DRAW12='1' OR DRAW13='1')) THEN
		R <= (OTHERS => '1');
		G <= (OTHERS => '0');
		B <= (OTHERS => '0');
		STOP <= '1';
	END IF;
	
	IF (HPOS < 1688) THEN
	HPOS <= HPOS + 1;
	ELSE
	HPOS <= 0;
		IF (VPOS < 1066) THEN
			VPOS <= VPOS + 1;
			ELSE
		
		IF(KEYS(0)='0')THEN
			START <= '1';
		END IF;
		
		IF(KEYS(1)='0')THEN
			START <= '1';
			STOP <= '0';
			PA_Y1 <= 0;
			PA_Y2 <= 0;
			PA_Y3 <= 0;
			PA_Y4 <= 0;
			PA_Y5 <= 0;
			PB_Y1 <= 1688; 
			PB_Y2 <= 1688; 
			PB_Y3 <= 1688; 
			PB_Y4 <= 1688; 
			PB_Y5 <= 1688; 
		END IF;
			
		IF(START='1' AND STOP='0')THEN
			IF(KEYS(0)='0')THEN
				SQ_Y1<=SQ_Y1 - 13;
			ELSE
				SQ_Y1<=SQ_Y1 + 8;
			END IF;
			
			PB_X1 <= PB_X1 - 6;
			PB_X2 <= PB_X2 - 6;
			PB_X3 <= PB_X3 - 6;
			PB_X4 <= PB_X4 - 6;
			PB_X5 <= PB_X5 - 6;
			PB_X6 <= PB_X6 - 6;
				
			PA_X1 <= PA_X1 - 6;
			PA_X2 <= PA_X2 - 6;
			PA_X3 <= PA_X3 - 6;
			PA_X4 <= PA_X4 - 6;
			PA_X5 <= PA_X5 - 6;
			PA_X6 <= PA_X6 - 6;
		END IF;
			--	END IF;
			-- IF(S(0)='1')THEN
				 
				 --IF(KEYS(1)='0')THEN
				 -- SQ_X1<=SQ_X1-5;
				-- END IF;
				 -- IF(KEYS(2)='0')THEN
				 -- SQ_Y1<=SQ_Y1-5;
				 --END IF;
				-- IF(KEYS(3)='0')THEN
				--  SQ_Y1<=SQ_Y1+5;
				-- END IF;  
			-- END IF;
			
			
			VPOS <= 0;
		END IF;
	END IF;
	
	IF (HPOS > 48 AND HPOS < 160) THEN
	HSYNC <= '0';
	ELSE
	HSYNC <= '1';
	END IF;
	
	IF (VPOS > 0 AND VPOS < 4) THEN
	VSYNC <= '0';
	ELSE
	VSYNC <= '1';
	END IF;
	
	IF ((HPOS > 0 AND HPOS < 408) OR (VPOS > 0 AND VPOS < 42)) THEN
	R <= (OTHERS=>'0');
	G <= (OTHERS=>'0');
	B <= (OTHERS=>'0');
	END IF;
	
END IF;
END PROCESS;
END MAIN;