library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

PACKAGE MY IS 
PROCEDURE SQ (
SIGNAL XCUR, YCUR, XPOS, YPOS: IN INTEGER;
SIGNAL RGB : OUT STD_LOGIC_VECTOR(3 downto 0);
SIGNAL DRAW: OUT STD_LOGIC
);
END MY

PACKAGE BODY MY IS
PROCEDURE SQ (
SIGNAL XCUR, YCUR, XPOS, YPOS: IN INTEGER;
SIGNAL RGB : OUT STD_LOGIC_VECTOR(3 downto 0);
SIGNAL DRAW: OUT STD_LOGIC) IS
BEGIN
IF (XCUR > XPOS AND XCUR < (XPOS + 100) AND YCUR > YPOS AND YCUR < (YPOS + 100)) THEN
RGB <= "1111";
DRAW <= '1';
ELSE
DRAW <= '0';
END IF;
END SQ;
END MY;